//----------------------+-------------------------------------------------------
// Filename             | compute_unit.sv
// File created on      | 09/02/2025
// Created by           | Sree Sankar E
//                      |
//                      |
//----------------------+-------------------------------------------------------
//
//------------------------------------------------------------------------------
// K Means Clustering Header
//------------------------------------------------------------------------------

`ifndef KMEANS_CLUSTER_H
`define KMEANS_CLUSTER_H

`endif